grammar edu:umn:cs:melt:exts:ableC:sed;

exports edu:umn:cs:melt:exts:ableC:sed:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:sed:concretesyntax;
